library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity rom is
  port
  (
    clk     : in std_logic;
    address : in unsigned(6 downto 0);
    data    : out unsigned(15 downto 0)
  );
end entity;
architecture rtl of rom is
  type mem is array (0 to 127) of unsigned(15 downto 0);
  constant rom_content : mem := (
        0 => "0110000000000010",
        1 => "0110000100000010",
        2 => "1011000000000000",
        3 => "0110000100000001",
        4 => "0001000000000000",
        5 => "1010000000000000",
        6 => "1011000000000000",
        7 => "0110000101111000",
        8 => "0101000000000000",
        9 => "1110111100100000",
        10 => "0110010000000000",
        11 => "0110001000000010",
        12 => "0110000100000010",
        13 => "0001001000000000",
        14 => "1010001000000000",
        15 => "1010010100000000",
        16 => "1011001000000000",
        17 => "0110000101111000",
        18 => "0101001000000000",
        19 => "1110111100000000",
        20 => "0110010000000000",
        21 => "0110001000000011",
        22 => "0110000100000011",
        23 => "0001001000000000",
        24 => "1010001000000000",
        25 => "1010010100000000",
        26 => "1011001000000000",
        27 => "0110000101111000",
        28 => "0101001000000000",
        29 => "1110111100000000",
        30 => "0110010000000000",
        31 => "0110001000000101",
        32 => "0110000100000101",
        33 => "0001001000000000",
        34 => "1010001000000000",
        35 => "1010010100000000",
        36 => "1011001000000000",
        37 => "0110000101111000",
        38 => "0101001000000000",
        39 => "1110111100000000",
        40 => "0110010000000000",
        41 => "0110001000000111",
        42 => "0110000100000111",
        43 => "0001001000000000",
        44 => "1010001000000000",
        45 => "1010010100000000",
        46 => "1011001000000000",
        47 => "0110000101111000",
        48 => "0101001000000000",
        49 => "1110111100000000",
        50 => "0110010000000000",
        51 => "0110001000001011",
        52 => "0110000100001011",
        53 => "0001001000000000",
        54 => "1010001000000000",
        55 => "1010010100000000",
        56 => "1011001000000000",
        57 => "0110000101111000",
        58 => "0101001000000000",
        59 => "1110111100000000",
        60 => "0110000000000001",
        61 => "0110000100000001",
        62 => "0001000000000000",
        63 => "1010000000000000",
        64 => "0111000000000000",
        65 => "1010111000000000",
        66 => "0110000101111000",
        67 => "0101000000000000",
        68 => "1110111100000000",
        others => (others => '0')
  );
begin
  process (clk)
  begin
    if (rising_edge(clk)) then
      data <= rom_content(to_integer(address));
    end if;
  end process;
end architecture;
