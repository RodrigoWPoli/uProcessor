library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity rom is
  port
  (
    clk     : in std_logic;
    address : in unsigned(6 downto 0);
    data    : out unsigned(15 downto 0)
  );
end entity;
architecture rtl of rom is
  type mem is array (0 to 127) of unsigned(15 downto 0);
  constant rom_content : mem := (
        0 => "0110000000000011",
        1 => "0110001000000111",
        2 => "0110010000001101",
        3 => "0110011000010000",
        4 => "0110100000011100",
        5 => "0110101000101000",
        6 => "0110110001100100",
        7 => "0110111001101110",
        8 => "0110000100100101",
        9 => "1011001000000000",
        10 => "0110000101011110",
        11 => "1011001000000000",
        12 => "0110000110111101",
        13 => "1011010000000000",
        14 => "0111000000000000",
        15 => "1010100000000000",
        16 => "0111101000000000",
        17 => "1010110000000000",
        18 => "0111000000000000",
        19 => "1010001000000000",
        20 => "0110000110100000",
        21 => "1011101000000000",
        22 => "0111001000000000",
        23 => "1010000000000000",
        24 => "0111011000000000",
        25 => "1010010000000000",
        26 => "0110000101100110",
        27 => "1011001000000000",
        28 => "0110000111110001",
        29 => "1011111000000000",
        30 => "0110000111001001",
        31 => "1011111000000000",
        32 => "0110000110111111",
        33 => "1011101000000000",
        34 => "0110000100010111",
        35 => "1011001000000000",
        36 => "0110000110000101",
        37 => "1011001000000000",
        38 => "0110000111110101",
        39 => "1011001000000000",
        40 => "0111001000000000",
        41 => "1010000000000000",
        42 => "0110000111110010",
        43 => "1011110000000000",
        44 => "0110000101011011",
        45 => "1011100000000000",
        46 => "0110000101000001",
        47 => "1011111000000000",
        48 => "0111100000000000",
        49 => "1010101000000000",
        50 => "0110000110100011",
        51 => "1011011000000000",
        52 => "0110000111010110",
        53 => "1011000000000000",
        54 => "0110000101101101",
        55 => "1011110000000000",
        56 => "0111111000000000",
        57 => "1010000000000000",
        58 => "0111011000000000",
        59 => "1010100000000000",
        60 => "0110000111111001",
        61 => "1011000000000000",
        62 => "0110000110000010",
        63 => "1011101000000000",
        64 => "0111001000000000",
        65 => "1010100000000000",
        66 => "0110000110011011",
        67 => "1011111000000000",
        68 => "0110000111000010",
        69 => "1011010000000000",
        70 => "0110000110110100",
        71 => "1011100000000000",
        72 => "0111000000000000",
        73 => "1010011000000000",
        74 => "0111100000000000",
        75 => "1010000000000000",
        76 => "0111110000000000",
        77 => "1010111000000000",
        78 => "0110000101010011",
        79 => "1011010000000000",
        80 => "0111010000000000",
        81 => "1010100000000000",
        82 => "0111101000000000",
        83 => "1010000000000000",
        84 => "0110000111100110",
        85 => "1011101000000000",
        86 => "0111010000000000",
        87 => "1010001000000000",
        88 => "0111010000000000",
        89 => "1010101000000000",
        90 => "0111111000000000",
        91 => "1010101000000000",
        92 => "0110000110110101",
        93 => "1011111000000000",
        94 => "0110000101110100",
        95 => "1011111000000000",
        96 => "0111110000000000",
        97 => "1010011000000000",
        98 => "0110000100111110",
        99 => "1011111000000000",
        100 => "0111111000000000",
        101 => "1010110000000000",
        102 => "0110000111111000",
        103 => "1011111000000000",
        104 => "0111111000000000",
        105 => "1010101000000000",
        106 => "0110000101100111",
        107 => "1011001000000000",
        others => (others => '0')
  );
begin
  process (clk)
  begin
    if (rising_edge(clk)) then
      data <= rom_content(to_integer(address));
    end if;
  end process;
end architecture;
