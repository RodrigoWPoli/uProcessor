library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity rom is
  port
  (
    clk     : in std_logic;
    address : in unsigned(6 downto 0);
    data    : out unsigned(15 downto 0)
  );
end entity;
architecture rtl of rom is
  type mem is array (0 to 127) of unsigned(15 downto 0);
  constant rom_content : mem := (
        0 => "0110000000000010", --ld, r0, 2
        1 => "0110000100000010", --ld, a, 2
        2 => "1011000000000000", --sw, r0
        3 => "0110000100000001", --ld, a, 1
        4 => "0001000000000000", --add, r0
        5 => "1010000000000000", --mov, r0
        6 => "1011000000000000", --sw, r0
        7 => "0110000101111000", --ld, a, 120
        8 => "0101000000000000", --cmp, r0
        9 => "1110111100100000", --blt, -7
        10 => "0110010000000000", --ld, r2, 0
        11 => "0110001000000010", --ld, r1, 2
        12 => "0110000100000010", --ld, a, 2
        13 => "0001001000000000", --add, r1
        14 => "1010001000000000", --mov, r1
        15 => "1010010100000000", --mov, a, r2
        16 => "1011001000000000", --sw, r1
        17 => "0110000101111000", --ld, a, 120
        18 => "0101001000000000", --cmp, r1
        19 => "1110111100000000", --blt, -8
        20 => "0110010000000000", --ld, r2, 0
        21 => "0110001000000011", --ld, r1, 3
        22 => "0110000100000011", --ld, a, 3
        23 => "0001001000000000", --add, r1
        24 => "1010001000000000", --mov, r1
        25 => "1010010100000000", --mov, a, r2
        26 => "1011001000000000", --sw, r1
        27 => "0110000101111000", --ld, a, 120
        28 => "0101001000000000", --cmp, r1
        29 => "1110111100000000", --blt, -8
        30 => "0110010000000000", --ld, r2, 0
        31 => "0110001000000101", --ld, r1, 5
        32 => "0110000100000101", --ld, a, 5
        33 => "0001001000000000", --add, r1
        34 => "1010001000000000", --mov, r1
        35 => "1010010100000000", --mov, a, r2
        36 => "1011001000000000", --sw, r1
        37 => "0110000101111000", --ld, a, 120
        38 => "0101001000000000", --cmp, r1
        39 => "1110111100000000", --blt, -8
        40 => "0110010000000000", --ld, r2, 0
        41 => "0110001000000111", --ld, r1, 7
        42 => "0110000100000111", --ld, a, 7
        43 => "0001001000000000", --add, r1
        44 => "1010001000000000", --mov, r1
        45 => "1010010100000000", --mov, a, r2
        46 => "1011001000000000", --sw, r1
        47 => "0110000101111000", --ld, a, 120
        48 => "0101001000000000", --cmp, r1
        49 => "1110111100000000", --blt, -8
        50 => "0110010000000000", --ld, r2, 0
        51 => "0110001000001011", --ld, r1, 11
        52 => "0110000100001011", --ld, a, 11
        53 => "0001001000000000", --add, r1
        54 => "1010001000000000", --mov, r1
        55 => "1010010100000000", --mov, a, r2
        56 => "1011001000000000", --sw, r1
        57 => "0110000101111000", --ld, a, 120
        58 => "0101001000000000", --cmp, r1
        59 => "1110111100000000", --blt, -8
        60 => "0110000000000001", --ld, r0, 1
        61 => "0110000100000001", --ld, a, 1
        62 => "0001000000000000", --add, r0
        63 => "1010000000000000", --mov, r0
        64 => "0111000000000000", --lw r0
        65 => "1010111000000000", --mov, r7
        66 => "0110000101111000", --ld, a, 120
        67 => "0101000000000000", --cmp, r0
        68 => "1110111100000000", --blt, -8
        others => (others => '0')
  );
begin
  process (clk)
  begin
    if (rising_edge(clk)) then
      data <= rom_content(to_integer(address));
    end if;
  end process;
end architecture;
